��l i b r a r y   i e e e   ;  
         u s e   i e e e . s t d _ l o g i c _ 1 1 6 4 . a l l   ;  
  
 e n t i t y   s e c o n d   i s  
     p o r t   ( )   ;  
 e n d   s e c o n d   ;    
  
 a r c h i t e c t u r e   a r c h   o f   s e c o n d   i s  
  
 b e g i n  
  
 e n d   a r c h i t e c t u r e   ;  
 